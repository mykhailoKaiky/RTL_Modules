library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity sinus_ROM is
Generic(length_ROM : natural; N_ROM_SIN : natural; N : natural);
Port ( 
        clk : in std_logic;
        reset : in std_logic;
        addr : in std_logic_vector(N_ROM_SIN-1 downto 0);
        output_ROM_data : out signed(N-1 downto 0) := (others => '0')
);
end sinus_ROM;

architecture Behavioral of sinus_ROM is
type SIN_ROM is array (0 to length_ROM-1) of signed(N-1 downto 0);

constant ROM : SIN_ROM :=
(
TO_SIGNED(    0,N),
TO_SIGNED(   50,N),
TO_SIGNED(  101,N),
TO_SIGNED(  151,N),
TO_SIGNED(  201,N),
TO_SIGNED(  251,N),
TO_SIGNED(  302,N),
TO_SIGNED(  352,N),
TO_SIGNED(  402,N),
TO_SIGNED(  452,N),
TO_SIGNED(  503,N),
TO_SIGNED(  553,N),
TO_SIGNED(  603,N),
TO_SIGNED(  653,N),
TO_SIGNED(  704,N),
TO_SIGNED(  754,N),
TO_SIGNED(  804,N),
TO_SIGNED(  854,N),
TO_SIGNED(  905,N),
TO_SIGNED(  955,N),
TO_SIGNED( 1005,N),
TO_SIGNED( 1055,N),
TO_SIGNED( 1106,N),
TO_SIGNED( 1156,N),
TO_SIGNED( 1206,N),
TO_SIGNED( 1256,N),
TO_SIGNED( 1307,N),
TO_SIGNED( 1357,N),
TO_SIGNED( 1407,N),
TO_SIGNED( 1457,N),
TO_SIGNED( 1507,N),
TO_SIGNED( 1558,N),
TO_SIGNED( 1608,N),
TO_SIGNED( 1658,N),
TO_SIGNED( 1708,N),
TO_SIGNED( 1758,N),
TO_SIGNED( 1809,N),
TO_SIGNED( 1859,N),
TO_SIGNED( 1909,N),
TO_SIGNED( 1959,N),
TO_SIGNED( 2009,N),
TO_SIGNED( 2060,N),
TO_SIGNED( 2110,N),
TO_SIGNED( 2160,N),
TO_SIGNED( 2210,N),
TO_SIGNED( 2260,N),
TO_SIGNED( 2310,N),
TO_SIGNED( 2360,N),
TO_SIGNED( 2411,N),
TO_SIGNED( 2461,N),
TO_SIGNED( 2511,N),
TO_SIGNED( 2561,N),
TO_SIGNED( 2611,N),
TO_SIGNED( 2661,N),
TO_SIGNED( 2711,N),
TO_SIGNED( 2761,N),
TO_SIGNED( 2811,N),
TO_SIGNED( 2861,N),
TO_SIGNED( 2912,N),
TO_SIGNED( 2962,N),
TO_SIGNED( 3012,N),
TO_SIGNED( 3062,N),
TO_SIGNED( 3112,N),
TO_SIGNED( 3162,N),
TO_SIGNED( 3212,N),
TO_SIGNED( 3262,N),
TO_SIGNED( 3312,N),
TO_SIGNED( 3362,N),
TO_SIGNED( 3412,N),
TO_SIGNED( 3462,N),
TO_SIGNED( 3512,N),
TO_SIGNED( 3562,N),
TO_SIGNED( 3612,N),
TO_SIGNED( 3662,N),
TO_SIGNED( 3712,N),
TO_SIGNED( 3762,N),
TO_SIGNED( 3812,N),
TO_SIGNED( 3861,N),
TO_SIGNED( 3911,N),
TO_SIGNED( 3961,N),
TO_SIGNED( 4011,N),
TO_SIGNED( 4061,N),
TO_SIGNED( 4111,N),
TO_SIGNED( 4161,N),
TO_SIGNED( 4211,N),
TO_SIGNED( 4260,N),
TO_SIGNED( 4310,N),
TO_SIGNED( 4360,N),
TO_SIGNED( 4410,N),
TO_SIGNED( 4460,N),
TO_SIGNED( 4510,N),
TO_SIGNED( 4559,N),
TO_SIGNED( 4609,N),
TO_SIGNED( 4659,N),
TO_SIGNED( 4709,N),
TO_SIGNED( 4758,N),
TO_SIGNED( 4808,N),
TO_SIGNED( 4858,N),
TO_SIGNED( 4907,N),
TO_SIGNED( 4957,N),
TO_SIGNED( 5007,N),
TO_SIGNED( 5057,N),
TO_SIGNED( 5106,N),
TO_SIGNED( 5156,N),
TO_SIGNED( 5205,N),
TO_SIGNED( 5255,N),
TO_SIGNED( 5305,N),
TO_SIGNED( 5354,N),
TO_SIGNED( 5404,N),
TO_SIGNED( 5453,N),
TO_SIGNED( 5503,N),
TO_SIGNED( 5553,N),
TO_SIGNED( 5602,N),
TO_SIGNED( 5652,N),
TO_SIGNED( 5701,N),
TO_SIGNED( 5751,N),
TO_SIGNED( 5800,N),
TO_SIGNED( 5850,N),
TO_SIGNED( 5899,N),
TO_SIGNED( 5948,N),
TO_SIGNED( 5998,N),
TO_SIGNED( 6047,N),
TO_SIGNED( 6097,N),
TO_SIGNED( 6146,N),
TO_SIGNED( 6195,N),
TO_SIGNED( 6245,N),
TO_SIGNED( 6294,N),
TO_SIGNED( 6343,N),
TO_SIGNED( 6393,N),
TO_SIGNED( 6442,N),
TO_SIGNED( 6491,N),
TO_SIGNED( 6541,N),
TO_SIGNED( 6590,N),
TO_SIGNED( 6639,N),
TO_SIGNED( 6688,N),
TO_SIGNED( 6737,N),
TO_SIGNED( 6787,N),
TO_SIGNED( 6836,N),
TO_SIGNED( 6885,N),
TO_SIGNED( 6934,N),
TO_SIGNED( 6983,N),
TO_SIGNED( 7032,N),
TO_SIGNED( 7081,N),
TO_SIGNED( 7130,N),
TO_SIGNED( 7180,N),
TO_SIGNED( 7229,N),
TO_SIGNED( 7278,N),
TO_SIGNED( 7327,N),
TO_SIGNED( 7376,N),
TO_SIGNED( 7425,N),
TO_SIGNED( 7473,N),
TO_SIGNED( 7522,N),
TO_SIGNED( 7571,N),
TO_SIGNED( 7620,N),
TO_SIGNED( 7669,N),
TO_SIGNED( 7718,N),
TO_SIGNED( 7767,N),
TO_SIGNED( 7816,N),
TO_SIGNED( 7864,N),
TO_SIGNED( 7913,N),
TO_SIGNED( 7962,N),
TO_SIGNED( 8011,N),
TO_SIGNED( 8059,N),
TO_SIGNED( 8108,N),
TO_SIGNED( 8157,N),
TO_SIGNED( 8206,N),
TO_SIGNED( 8254,N),
TO_SIGNED( 8303,N),
TO_SIGNED( 8351,N),
TO_SIGNED( 8400,N),
TO_SIGNED( 8449,N),
TO_SIGNED( 8497,N),
TO_SIGNED( 8546,N),
TO_SIGNED( 8594,N),
TO_SIGNED( 8643,N),
TO_SIGNED( 8691,N),
TO_SIGNED( 8740,N),
TO_SIGNED( 8788,N),
TO_SIGNED( 8836,N),
TO_SIGNED( 8885,N),
TO_SIGNED( 8933,N),
TO_SIGNED( 8982,N),
TO_SIGNED( 9030,N),
TO_SIGNED( 9078,N),
TO_SIGNED( 9127,N),
TO_SIGNED( 9175,N),
TO_SIGNED( 9223,N),
TO_SIGNED( 9271,N),
TO_SIGNED( 9319,N),
TO_SIGNED( 9368,N),
TO_SIGNED( 9416,N),
TO_SIGNED( 9464,N),
TO_SIGNED( 9512,N),
TO_SIGNED( 9560,N),
TO_SIGNED( 9608,N),
TO_SIGNED( 9656,N),
TO_SIGNED( 9704,N),
TO_SIGNED( 9752,N),
TO_SIGNED( 9800,N),
TO_SIGNED( 9848,N),
TO_SIGNED( 9896,N),
TO_SIGNED( 9944,N),
TO_SIGNED( 9992,N),
TO_SIGNED(10040,N),
TO_SIGNED(10088,N),
TO_SIGNED(10135,N),
TO_SIGNED(10183,N),
TO_SIGNED(10231,N),
TO_SIGNED(10279,N),
TO_SIGNED(10326,N),
TO_SIGNED(10374,N),
TO_SIGNED(10422,N),
TO_SIGNED(10469,N),
TO_SIGNED(10517,N),
TO_SIGNED(10565,N),
TO_SIGNED(10612,N),
TO_SIGNED(10660,N),
TO_SIGNED(10707,N),
TO_SIGNED(10755,N),
TO_SIGNED(10802,N),
TO_SIGNED(10850,N),
TO_SIGNED(10897,N),
TO_SIGNED(10945,N),
TO_SIGNED(10992,N),
TO_SIGNED(11039,N),
TO_SIGNED(11087,N),
TO_SIGNED(11134,N),
TO_SIGNED(11181,N),
TO_SIGNED(11228,N),
TO_SIGNED(11276,N),
TO_SIGNED(11323,N),
TO_SIGNED(11370,N),
TO_SIGNED(11417,N),
TO_SIGNED(11464,N),
TO_SIGNED(11511,N),
TO_SIGNED(11558,N),
TO_SIGNED(11605,N),
TO_SIGNED(11652,N),
TO_SIGNED(11699,N),
TO_SIGNED(11746,N),
TO_SIGNED(11793,N),
TO_SIGNED(11840,N),
TO_SIGNED(11887,N),
TO_SIGNED(11934,N),
TO_SIGNED(11980,N),
TO_SIGNED(12027,N),
TO_SIGNED(12074,N),
TO_SIGNED(12121,N),
TO_SIGNED(12167,N),
TO_SIGNED(12214,N),
TO_SIGNED(12261,N),
TO_SIGNED(12307,N),
TO_SIGNED(12354,N),
TO_SIGNED(12400,N),
TO_SIGNED(12447,N),
TO_SIGNED(12493,N),
TO_SIGNED(12540,N),
TO_SIGNED(12586,N),
TO_SIGNED(12633,N),
TO_SIGNED(12679,N),
TO_SIGNED(12725,N),
TO_SIGNED(12772,N),
TO_SIGNED(12818,N),
TO_SIGNED(12864,N),
TO_SIGNED(12910,N),
TO_SIGNED(12957,N),
TO_SIGNED(13003,N),
TO_SIGNED(13049,N),
TO_SIGNED(13095,N),
TO_SIGNED(13141,N),
TO_SIGNED(13187,N),
TO_SIGNED(13233,N),
TO_SIGNED(13279,N),
TO_SIGNED(13325,N),
TO_SIGNED(13371,N),
TO_SIGNED(13417,N),
TO_SIGNED(13463,N),
TO_SIGNED(13508,N),
TO_SIGNED(13554,N),
TO_SIGNED(13600,N),
TO_SIGNED(13646,N),
TO_SIGNED(13691,N),
TO_SIGNED(13737,N),
TO_SIGNED(13783,N),
TO_SIGNED(13828,N),
TO_SIGNED(13874,N),
TO_SIGNED(13919,N),
TO_SIGNED(13965,N),
TO_SIGNED(14010,N),
TO_SIGNED(14056,N),
TO_SIGNED(14101,N),
TO_SIGNED(14146,N),
TO_SIGNED(14192,N),
TO_SIGNED(14237,N),
TO_SIGNED(14282,N),
TO_SIGNED(14327,N),
TO_SIGNED(14373,N),
TO_SIGNED(14418,N),
TO_SIGNED(14463,N),
TO_SIGNED(14508,N),
TO_SIGNED(14553,N),
TO_SIGNED(14598,N),
TO_SIGNED(14643,N),
TO_SIGNED(14688,N),
TO_SIGNED(14733,N),
TO_SIGNED(14778,N),
TO_SIGNED(14823,N),
TO_SIGNED(14867,N),
TO_SIGNED(14912,N),
TO_SIGNED(14957,N),
TO_SIGNED(15002,N),
TO_SIGNED(15046,N),
TO_SIGNED(15091,N),
TO_SIGNED(15136,N),
TO_SIGNED(15180,N),
TO_SIGNED(15225,N),
TO_SIGNED(15269,N),
TO_SIGNED(15314,N),
TO_SIGNED(15358,N),
TO_SIGNED(15402,N),
TO_SIGNED(15447,N),
TO_SIGNED(15491,N),
TO_SIGNED(15535,N),
TO_SIGNED(15580,N),
TO_SIGNED(15624,N),
TO_SIGNED(15668,N),
TO_SIGNED(15712,N),
TO_SIGNED(15756,N),
TO_SIGNED(15800,N),
TO_SIGNED(15844,N),
TO_SIGNED(15888,N),
TO_SIGNED(15932,N),
TO_SIGNED(15976,N),
TO_SIGNED(16020,N),
TO_SIGNED(16064,N),
TO_SIGNED(16108,N),
TO_SIGNED(16151,N),
TO_SIGNED(16195,N),
TO_SIGNED(16239,N),
TO_SIGNED(16282,N),
TO_SIGNED(16326,N),
TO_SIGNED(16369,N),
TO_SIGNED(16413,N),
TO_SIGNED(16456,N),
TO_SIGNED(16500,N),
TO_SIGNED(16543,N),
TO_SIGNED(16587,N),
TO_SIGNED(16630,N),
TO_SIGNED(16673,N),
TO_SIGNED(16717,N),
TO_SIGNED(16760,N),
TO_SIGNED(16803,N),
TO_SIGNED(16846,N),
TO_SIGNED(16889,N),
TO_SIGNED(16932,N),
TO_SIGNED(16975,N),
TO_SIGNED(17018,N),
TO_SIGNED(17061,N),
TO_SIGNED(17104,N),
TO_SIGNED(17147,N),
TO_SIGNED(17190,N),
TO_SIGNED(17233,N),
TO_SIGNED(17275,N),
TO_SIGNED(17318,N),
TO_SIGNED(17361,N),
TO_SIGNED(17403,N),
TO_SIGNED(17446,N),
TO_SIGNED(17488,N),
TO_SIGNED(17531,N),
TO_SIGNED(17573,N),
TO_SIGNED(17616,N),
TO_SIGNED(17658,N),
TO_SIGNED(17700,N),
TO_SIGNED(17743,N),
TO_SIGNED(17785,N),
TO_SIGNED(17827,N),
TO_SIGNED(17869,N),
TO_SIGNED(17911,N),
TO_SIGNED(17953,N),
TO_SIGNED(17995,N),
TO_SIGNED(18037,N),
TO_SIGNED(18079,N),
TO_SIGNED(18121,N),
TO_SIGNED(18163,N),
TO_SIGNED(18205,N),
TO_SIGNED(18247,N),
TO_SIGNED(18288,N),
TO_SIGNED(18330,N),
TO_SIGNED(18372,N),
TO_SIGNED(18413,N),
TO_SIGNED(18455,N),
TO_SIGNED(18496,N),
TO_SIGNED(18538,N),
TO_SIGNED(18579,N),
TO_SIGNED(18621,N),
TO_SIGNED(18662,N),
TO_SIGNED(18703,N),
TO_SIGNED(18745,N),
TO_SIGNED(18786,N),
TO_SIGNED(18827,N),
TO_SIGNED(18868,N),
TO_SIGNED(18909,N),
TO_SIGNED(18950,N),
TO_SIGNED(18991,N),
TO_SIGNED(19032,N),
TO_SIGNED(19073,N),
TO_SIGNED(19114,N),
TO_SIGNED(19155,N),
TO_SIGNED(19195,N),
TO_SIGNED(19236,N),
TO_SIGNED(19277,N),
TO_SIGNED(19317,N),
TO_SIGNED(19358,N),
TO_SIGNED(19399,N),
TO_SIGNED(19439,N),
TO_SIGNED(19479,N),
TO_SIGNED(19520,N),
TO_SIGNED(19560,N),
TO_SIGNED(19601,N),
TO_SIGNED(19641,N),
TO_SIGNED(19681,N),
TO_SIGNED(19721,N),
TO_SIGNED(19761,N),
TO_SIGNED(19801,N),
TO_SIGNED(19841,N),
TO_SIGNED(19881,N),
TO_SIGNED(19921,N),
TO_SIGNED(19961,N),
TO_SIGNED(20001,N),
TO_SIGNED(20041,N),
TO_SIGNED(20081,N),
TO_SIGNED(20120,N),
TO_SIGNED(20160,N),
TO_SIGNED(20200,N),
TO_SIGNED(20239,N),
TO_SIGNED(20279,N),
TO_SIGNED(20318,N),
TO_SIGNED(20357,N),
TO_SIGNED(20397,N),
TO_SIGNED(20436,N),
TO_SIGNED(20475,N),
TO_SIGNED(20515,N),
TO_SIGNED(20554,N),
TO_SIGNED(20593,N),
TO_SIGNED(20632,N),
TO_SIGNED(20671,N),
TO_SIGNED(20710,N),
TO_SIGNED(20749,N),
TO_SIGNED(20788,N),
TO_SIGNED(20827,N),
TO_SIGNED(20865,N),
TO_SIGNED(20904,N),
TO_SIGNED(20943,N),
TO_SIGNED(20981,N),
TO_SIGNED(21020,N),
TO_SIGNED(21059,N),
TO_SIGNED(21097,N),
TO_SIGNED(21136,N),
TO_SIGNED(21174,N),
TO_SIGNED(21212,N),
TO_SIGNED(21251,N),
TO_SIGNED(21289,N),
TO_SIGNED(21327,N),
TO_SIGNED(21365,N),
TO_SIGNED(21403,N),
TO_SIGNED(21441,N),
TO_SIGNED(21479,N),
TO_SIGNED(21517,N),
TO_SIGNED(21555,N),
TO_SIGNED(21593,N),
TO_SIGNED(21631,N),
TO_SIGNED(21668,N),
TO_SIGNED(21706,N),
TO_SIGNED(21744,N),
TO_SIGNED(21781,N),
TO_SIGNED(21819,N),
TO_SIGNED(21856,N),
TO_SIGNED(21894,N),
TO_SIGNED(21931,N),
TO_SIGNED(21968,N),
TO_SIGNED(22006,N),
TO_SIGNED(22043,N),
TO_SIGNED(22080,N),
TO_SIGNED(22117,N),
TO_SIGNED(22154,N),
TO_SIGNED(22191,N),
TO_SIGNED(22228,N),
TO_SIGNED(22265,N),
TO_SIGNED(22302,N),
TO_SIGNED(22339,N),
TO_SIGNED(22375,N),
TO_SIGNED(22412,N),
TO_SIGNED(22449,N),
TO_SIGNED(22485,N),
TO_SIGNED(22522,N),
TO_SIGNED(22558,N),
TO_SIGNED(22595,N),
TO_SIGNED(22631,N),
TO_SIGNED(22668,N),
TO_SIGNED(22704,N),
TO_SIGNED(22740,N),
TO_SIGNED(22776,N),
TO_SIGNED(22812,N),
TO_SIGNED(22848,N),
TO_SIGNED(22884,N),
TO_SIGNED(22920,N),
TO_SIGNED(22956,N),
TO_SIGNED(22992,N),
TO_SIGNED(23028,N),
TO_SIGNED(23064,N),
TO_SIGNED(23099,N),
TO_SIGNED(23135,N),
TO_SIGNED(23170,N),
TO_SIGNED(23206,N),
TO_SIGNED(23241,N),
TO_SIGNED(23277,N),
TO_SIGNED(23312,N),
TO_SIGNED(23348,N),
TO_SIGNED(23383,N),
TO_SIGNED(23418,N),
TO_SIGNED(23453,N),
TO_SIGNED(23488,N),
TO_SIGNED(23523,N),
TO_SIGNED(23558,N),
TO_SIGNED(23593,N),
TO_SIGNED(23628,N),
TO_SIGNED(23663,N),
TO_SIGNED(23697,N),
TO_SIGNED(23732,N),
TO_SIGNED(23767,N),
TO_SIGNED(23801,N),
TO_SIGNED(23836,N),
TO_SIGNED(23870,N),
TO_SIGNED(23905,N),
TO_SIGNED(23939,N),
TO_SIGNED(23973,N),
TO_SIGNED(24008,N),
TO_SIGNED(24042,N),
TO_SIGNED(24076,N),
TO_SIGNED(24110,N),
TO_SIGNED(24144,N),
TO_SIGNED(24178,N),
TO_SIGNED(24212,N),
TO_SIGNED(24246,N),
TO_SIGNED(24279,N),
TO_SIGNED(24313,N),
TO_SIGNED(24347,N),
TO_SIGNED(24380,N),
TO_SIGNED(24414,N),
TO_SIGNED(24448,N),
TO_SIGNED(24481,N),
TO_SIGNED(24514,N),
TO_SIGNED(24548,N),
TO_SIGNED(24581,N),
TO_SIGNED(24614,N),
TO_SIGNED(24647,N),
TO_SIGNED(24680,N),
TO_SIGNED(24713,N),
TO_SIGNED(24746,N),
TO_SIGNED(24779,N),
TO_SIGNED(24812,N),
TO_SIGNED(24845,N),
TO_SIGNED(24878,N),
TO_SIGNED(24910,N),
TO_SIGNED(24943,N),
TO_SIGNED(24976,N),
TO_SIGNED(25008,N),
TO_SIGNED(25041,N),
TO_SIGNED(25073,N),
TO_SIGNED(25105,N),
TO_SIGNED(25138,N),
TO_SIGNED(25170,N),
TO_SIGNED(25202,N),
TO_SIGNED(25234,N),
TO_SIGNED(25266,N),
TO_SIGNED(25298,N),
TO_SIGNED(25330,N),
TO_SIGNED(25362,N),
TO_SIGNED(25394,N),
TO_SIGNED(25425,N),
TO_SIGNED(25457,N),
TO_SIGNED(25489,N),
TO_SIGNED(25520,N),
TO_SIGNED(25552,N),
TO_SIGNED(25583,N),
TO_SIGNED(25615,N),
TO_SIGNED(25646,N),
TO_SIGNED(25677,N),
TO_SIGNED(25708,N),
TO_SIGNED(25739,N),
TO_SIGNED(25771,N),
TO_SIGNED(25802,N),
TO_SIGNED(25833,N),
TO_SIGNED(25863,N),
TO_SIGNED(25894,N),
TO_SIGNED(25925,N),
TO_SIGNED(25956,N),
TO_SIGNED(25986,N),
TO_SIGNED(26017,N),
TO_SIGNED(26048,N),
TO_SIGNED(26078,N),
TO_SIGNED(26108,N),
TO_SIGNED(26139,N),
TO_SIGNED(26169,N),
TO_SIGNED(26199,N),
TO_SIGNED(26229,N),
TO_SIGNED(26259,N),
TO_SIGNED(26290,N),
TO_SIGNED(26320,N),
TO_SIGNED(26349,N),
TO_SIGNED(26379,N),
TO_SIGNED(26409,N),
TO_SIGNED(26439,N),
TO_SIGNED(26468,N),
TO_SIGNED(26498,N),
TO_SIGNED(26528,N),
TO_SIGNED(26557,N),
TO_SIGNED(26586,N),
TO_SIGNED(26616,N),
TO_SIGNED(26645,N),
TO_SIGNED(26674,N),
TO_SIGNED(26704,N),
TO_SIGNED(26733,N),
TO_SIGNED(26762,N),
TO_SIGNED(26791,N),
TO_SIGNED(26820,N),
TO_SIGNED(26848,N),
TO_SIGNED(26877,N),
TO_SIGNED(26906,N),
TO_SIGNED(26935,N),
TO_SIGNED(26963,N),
TO_SIGNED(26992,N),
TO_SIGNED(27020,N),
TO_SIGNED(27049,N),
TO_SIGNED(27077,N),
TO_SIGNED(27105,N),
TO_SIGNED(27133,N),
TO_SIGNED(27162,N),
TO_SIGNED(27190,N),
TO_SIGNED(27218,N),
TO_SIGNED(27246,N),
TO_SIGNED(27273,N),
TO_SIGNED(27301,N),
TO_SIGNED(27329,N),
TO_SIGNED(27357,N),
TO_SIGNED(27384,N),
TO_SIGNED(27412,N),
TO_SIGNED(27440,N),
TO_SIGNED(27467,N),
TO_SIGNED(27494,N),
TO_SIGNED(27522,N),
TO_SIGNED(27549,N),
TO_SIGNED(27576,N),
TO_SIGNED(27603,N),
TO_SIGNED(27630,N),
TO_SIGNED(27657,N),
TO_SIGNED(27684,N),
TO_SIGNED(27711,N),
TO_SIGNED(27738,N),
TO_SIGNED(27765,N),
TO_SIGNED(27791,N),
TO_SIGNED(27818,N),
TO_SIGNED(27844,N),
TO_SIGNED(27871,N),
TO_SIGNED(27897,N),
TO_SIGNED(27924,N),
TO_SIGNED(27950,N),
TO_SIGNED(27976,N),
TO_SIGNED(28002,N),
TO_SIGNED(28028,N),
TO_SIGNED(28054,N),
TO_SIGNED(28080,N),
TO_SIGNED(28106,N),
TO_SIGNED(28132,N),
TO_SIGNED(28158,N),
TO_SIGNED(28183,N),
TO_SIGNED(28209,N),
TO_SIGNED(28234,N),
TO_SIGNED(28260,N),
TO_SIGNED(28285,N),
TO_SIGNED(28311,N),
TO_SIGNED(28336,N),
TO_SIGNED(28361,N),
TO_SIGNED(28386,N),
TO_SIGNED(28411,N),
TO_SIGNED(28436,N),
TO_SIGNED(28461,N),
TO_SIGNED(28486,N),
TO_SIGNED(28511,N),
TO_SIGNED(28536,N),
TO_SIGNED(28560,N),
TO_SIGNED(28585,N),
TO_SIGNED(28610,N),
TO_SIGNED(28634,N),
TO_SIGNED(28658,N),
TO_SIGNED(28683,N),
TO_SIGNED(28707,N),
TO_SIGNED(28731,N),
TO_SIGNED(28755,N),
TO_SIGNED(28779,N),
TO_SIGNED(28803,N),
TO_SIGNED(28827,N),
TO_SIGNED(28851,N),
TO_SIGNED(28875,N),
TO_SIGNED(28899,N),
TO_SIGNED(28922,N),
TO_SIGNED(28946,N),
TO_SIGNED(28970,N),
TO_SIGNED(28993,N),
TO_SIGNED(29016,N),
TO_SIGNED(29040,N),
TO_SIGNED(29063,N),
TO_SIGNED(29086,N),
TO_SIGNED(29109,N),
TO_SIGNED(29132,N),
TO_SIGNED(29155,N),
TO_SIGNED(29178,N),
TO_SIGNED(29201,N),
TO_SIGNED(29224,N),
TO_SIGNED(29247,N),
TO_SIGNED(29269,N),
TO_SIGNED(29292,N),
TO_SIGNED(29314,N),
TO_SIGNED(29337,N),
TO_SIGNED(29359,N),
TO_SIGNED(29381,N),
TO_SIGNED(29404,N),
TO_SIGNED(29426,N),
TO_SIGNED(29448,N),
TO_SIGNED(29470,N),
TO_SIGNED(29492,N),
TO_SIGNED(29514,N),
TO_SIGNED(29535,N),
TO_SIGNED(29557,N),
TO_SIGNED(29579,N),
TO_SIGNED(29600,N),
TO_SIGNED(29622,N),
TO_SIGNED(29643,N),
TO_SIGNED(29665,N),
TO_SIGNED(29686,N),
TO_SIGNED(29707,N),
TO_SIGNED(29729,N),
TO_SIGNED(29750,N),
TO_SIGNED(29771,N),
TO_SIGNED(29792,N),
TO_SIGNED(29813,N),
TO_SIGNED(29833,N),
TO_SIGNED(29854,N),
TO_SIGNED(29875,N),
TO_SIGNED(29895,N),
TO_SIGNED(29916,N),
TO_SIGNED(29936,N),
TO_SIGNED(29957,N),
TO_SIGNED(29977,N),
TO_SIGNED(29997,N),
TO_SIGNED(30018,N),
TO_SIGNED(30038,N),
TO_SIGNED(30058,N),
TO_SIGNED(30078,N),
TO_SIGNED(30098,N),
TO_SIGNED(30118,N),
TO_SIGNED(30137,N),
TO_SIGNED(30157,N),
TO_SIGNED(30177,N),
TO_SIGNED(30196,N),
TO_SIGNED(30216,N),
TO_SIGNED(30235,N),
TO_SIGNED(30254,N),
TO_SIGNED(30274,N),
TO_SIGNED(30293,N),
TO_SIGNED(30312,N),
TO_SIGNED(30331,N),
TO_SIGNED(30350,N),
TO_SIGNED(30369,N),
TO_SIGNED(30388,N),
TO_SIGNED(30407,N),
TO_SIGNED(30425,N),
TO_SIGNED(30444,N),
TO_SIGNED(30462,N),
TO_SIGNED(30481,N),
TO_SIGNED(30499,N),
TO_SIGNED(30518,N),
TO_SIGNED(30536,N),
TO_SIGNED(30554,N),
TO_SIGNED(30572,N),
TO_SIGNED(30590,N),
TO_SIGNED(30608,N),
TO_SIGNED(30626,N),
TO_SIGNED(30644,N),
TO_SIGNED(30662,N),
TO_SIGNED(30680,N),
TO_SIGNED(30697,N),
TO_SIGNED(30715,N),
TO_SIGNED(30732,N),
TO_SIGNED(30750,N),
TO_SIGNED(30767,N),
TO_SIGNED(30784,N),
TO_SIGNED(30801,N),
TO_SIGNED(30819,N),
TO_SIGNED(30836,N),
TO_SIGNED(30853,N),
TO_SIGNED(30869,N),
TO_SIGNED(30886,N),
TO_SIGNED(30903,N),
TO_SIGNED(30920,N),
TO_SIGNED(30936,N),
TO_SIGNED(30953,N),
TO_SIGNED(30969,N),
TO_SIGNED(30986,N),
TO_SIGNED(31002,N),
TO_SIGNED(31018,N),
TO_SIGNED(31034,N),
TO_SIGNED(31050,N),
TO_SIGNED(31067,N),
TO_SIGNED(31082,N),
TO_SIGNED(31098,N),
TO_SIGNED(31114,N),
TO_SIGNED(31130,N),
TO_SIGNED(31146,N),
TO_SIGNED(31161,N),
TO_SIGNED(31177,N),
TO_SIGNED(31192,N),
TO_SIGNED(31207,N),
TO_SIGNED(31223,N),
TO_SIGNED(31238,N),
TO_SIGNED(31253,N),
TO_SIGNED(31268,N),
TO_SIGNED(31283,N),
TO_SIGNED(31298,N),
TO_SIGNED(31313,N),
TO_SIGNED(31328,N),
TO_SIGNED(31342,N),
TO_SIGNED(31357,N),
TO_SIGNED(31372,N),
TO_SIGNED(31386,N),
TO_SIGNED(31400,N),
TO_SIGNED(31415,N),
TO_SIGNED(31429,N),
TO_SIGNED(31443,N),
TO_SIGNED(31457,N),
TO_SIGNED(31471,N),
TO_SIGNED(31485,N),
TO_SIGNED(31499,N),
TO_SIGNED(31513,N),
TO_SIGNED(31527,N),
TO_SIGNED(31540,N),
TO_SIGNED(31554,N),
TO_SIGNED(31568,N),
TO_SIGNED(31581,N),
TO_SIGNED(31594,N),
TO_SIGNED(31608,N),
TO_SIGNED(31621,N),
TO_SIGNED(31634,N),
TO_SIGNED(31647,N),
TO_SIGNED(31660,N),
TO_SIGNED(31673,N),
TO_SIGNED(31686,N),
TO_SIGNED(31699,N),
TO_SIGNED(31711,N),
TO_SIGNED(31724,N),
TO_SIGNED(31737,N),
TO_SIGNED(31749,N),
TO_SIGNED(31761,N),
TO_SIGNED(31774,N),
TO_SIGNED(31786,N),
TO_SIGNED(31798,N),
TO_SIGNED(31810,N),
TO_SIGNED(31822,N),
TO_SIGNED(31834,N),
TO_SIGNED(31846,N),
TO_SIGNED(31858,N),
TO_SIGNED(31870,N),
TO_SIGNED(31881,N),
TO_SIGNED(31893,N),
TO_SIGNED(31904,N),
TO_SIGNED(31916,N),
TO_SIGNED(31927,N),
TO_SIGNED(31938,N),
TO_SIGNED(31950,N),
TO_SIGNED(31961,N),
TO_SIGNED(31972,N),
TO_SIGNED(31983,N),
TO_SIGNED(31994,N),
TO_SIGNED(32005,N),
TO_SIGNED(32015,N),
TO_SIGNED(32026,N),
TO_SIGNED(32037,N),
TO_SIGNED(32047,N),
TO_SIGNED(32058,N),
TO_SIGNED(32068,N),
TO_SIGNED(32078,N),
TO_SIGNED(32088,N),
TO_SIGNED(32099,N),
TO_SIGNED(32109,N),
TO_SIGNED(32119,N),
TO_SIGNED(32129,N),
TO_SIGNED(32138,N),
TO_SIGNED(32148,N),
TO_SIGNED(32158,N),
TO_SIGNED(32167,N),
TO_SIGNED(32177,N),
TO_SIGNED(32186,N),
TO_SIGNED(32196,N),
TO_SIGNED(32205,N),
TO_SIGNED(32214,N),
TO_SIGNED(32224,N),
TO_SIGNED(32233,N),
TO_SIGNED(32242,N),
TO_SIGNED(32251,N),
TO_SIGNED(32259,N),
TO_SIGNED(32268,N),
TO_SIGNED(32277,N),
TO_SIGNED(32286,N),
TO_SIGNED(32294,N),
TO_SIGNED(32303,N),
TO_SIGNED(32311,N),
TO_SIGNED(32319,N),
TO_SIGNED(32328,N),
TO_SIGNED(32336,N),
TO_SIGNED(32344,N),
TO_SIGNED(32352,N),
TO_SIGNED(32360,N),
TO_SIGNED(32368,N),
TO_SIGNED(32376,N),
TO_SIGNED(32383,N),
TO_SIGNED(32391,N),
TO_SIGNED(32398,N),
TO_SIGNED(32406,N),
TO_SIGNED(32413,N),
TO_SIGNED(32421,N),
TO_SIGNED(32428,N),
TO_SIGNED(32435,N),
TO_SIGNED(32442,N),
TO_SIGNED(32449,N),
TO_SIGNED(32456,N),
TO_SIGNED(32463,N),
TO_SIGNED(32470,N),
TO_SIGNED(32477,N),
TO_SIGNED(32483,N),
TO_SIGNED(32490,N),
TO_SIGNED(32496,N),
TO_SIGNED(32503,N),
TO_SIGNED(32509,N),
TO_SIGNED(32515,N),
TO_SIGNED(32522,N),
TO_SIGNED(32528,N),
TO_SIGNED(32534,N),
TO_SIGNED(32540,N),
TO_SIGNED(32546,N),
TO_SIGNED(32551,N),
TO_SIGNED(32557,N),
TO_SIGNED(32563,N),
TO_SIGNED(32568,N),
TO_SIGNED(32574,N),
TO_SIGNED(32579,N),
TO_SIGNED(32585,N),
TO_SIGNED(32590,N),
TO_SIGNED(32595,N),
TO_SIGNED(32600,N),
TO_SIGNED(32605,N),
TO_SIGNED(32610,N),
TO_SIGNED(32615,N),
TO_SIGNED(32620,N),
TO_SIGNED(32625,N),
TO_SIGNED(32629,N),
TO_SIGNED(32634,N),
TO_SIGNED(32638,N),
TO_SIGNED(32643,N),
TO_SIGNED(32647,N),
TO_SIGNED(32651,N),
TO_SIGNED(32656,N),
TO_SIGNED(32660,N),
TO_SIGNED(32664,N),
TO_SIGNED(32668,N),
TO_SIGNED(32672,N),
TO_SIGNED(32675,N),
TO_SIGNED(32679,N),
TO_SIGNED(32683,N),
TO_SIGNED(32686,N),
TO_SIGNED(32690,N),
TO_SIGNED(32693,N),
TO_SIGNED(32697,N),
TO_SIGNED(32700,N),
TO_SIGNED(32703,N),
TO_SIGNED(32706,N),
TO_SIGNED(32709,N),
TO_SIGNED(32712,N),
TO_SIGNED(32715,N),
TO_SIGNED(32718,N),
TO_SIGNED(32721,N),
TO_SIGNED(32723,N),
TO_SIGNED(32726,N),
TO_SIGNED(32729,N),
TO_SIGNED(32731,N),
TO_SIGNED(32733,N),
TO_SIGNED(32736,N),
TO_SIGNED(32738,N),
TO_SIGNED(32740,N),
TO_SIGNED(32742,N),
TO_SIGNED(32744,N),
TO_SIGNED(32746,N),
TO_SIGNED(32748,N),
TO_SIGNED(32749,N),
TO_SIGNED(32751,N),
TO_SIGNED(32753,N),
TO_SIGNED(32754,N),
TO_SIGNED(32756,N),
TO_SIGNED(32757,N),
TO_SIGNED(32758,N),
TO_SIGNED(32759,N),
TO_SIGNED(32760,N),
TO_SIGNED(32761,N),
TO_SIGNED(32762,N),
TO_SIGNED(32763,N),
TO_SIGNED(32764,N),
TO_SIGNED(32765,N),
TO_SIGNED(32766,N),
TO_SIGNED(32766,N),
TO_SIGNED(32767,N),
TO_SIGNED(32767,N),
TO_SIGNED(32767,N),
TO_SIGNED(32767,N),
TO_SIGNED(32767,N),
TO_SIGNED(32767,N)
);
begin
process(clk,reset)
begin
if reset = '1' then
     output_ROM_data <= (others => '0');
elsif rising_edge(clk) then
    output_ROM_data <= ROM(TO_INTEGER(UNSIGNED(addr)));
end if;
end process;

end Behavioral;
